package FIFO_shared_pkg;
	parameter FIFO_WIDTH=16;
	parameter FIFO_DEPTH=32;
endpackage